module core_module
(
    input [71:0]            data_i,

    output  [7:0]           pixel_o,
    output                  core_valid_i
);



endmodule