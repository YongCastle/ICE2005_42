`timescale 1ns / 1ps

module SOBER_TOP
(
    
);


endmodule