module vga_buffer
(
)

endmodule